// Title         : vending_machine_def.v
// Author      : Jae-Eon Jo (Jojaeeon@postech.ac.kr) 
//					Dongup Kwon (nankdu7@postech.ac.kr)

// Macro constants (prefix k & CamelCase)
`define kTotalBits 31
  
`define kItemBits 8
`define kNumItems 4

`define kCoinBits 8
`define kNumCoins 3

`define kWaitTime 100